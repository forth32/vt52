//************************************************************
//*   Текстовый видеоадаптер с VGA-выходом
//************************************************************
module vga (
// шина wishbone
   input						wb_clk_i,	// тактовая частота шины
	input						wb_rst_i,	// сброс
	input	 [15:0]			wb_adr_i,	// адрес 
	input	 [15:0]			wb_dat_i,	// входные данные
   output reg [15:0]		wb_dat_o,	// выходные данные
	input						wb_cyc_i,	// начало цикла шины
	input	  					wb_we_i,		// разрешение записи (0 - чтение)
	input						wb_stb_i,	// строб цикла шины
	input	 [1:0]	      wb_sel_i,   // выбор конкретных байтов для записи - старший, младший или оба
	output reg				wb_ack_o,	// подтверждение выбора устройства
   // VGA      
   output reg vga_hsync,         // строчный синхросингал
   output reg vga_vsync,         // кадровый синхросигнал 
   output vgar,             // видеовыход красный
   output vgag,             // видеовыход зеленый
   output vgab,             // видеовыход синий
   // управление
   input[12:0] cursor,           // адрес курсора
	input lmode,                  // 0 - 24 строки, 1 - 38 строк
	input cursor_on,              // 0 - курсор невидим, 1 - отображается
	input cursor_type,           // форма курсора, 0 - подчеркивание, 1 - блок
   input flash,                 // импульсы переключения видимости мерцающих символов
	
   input clk50mhz                // тактовый сигнал 50 Мгц
);

	// двухпортовый видеобуфер
   reg[7:0] vram_even[0:2047]; 			// четные байты
   reg[7:0] vram_odd[0:2047]; 			// нечетные байты
	
   reg vgaclk;                // пиксельный синхросигнал (тактовая частота видеовыхода)
   reg[10:0] col;             // текущий столбец
   reg[9:0] row;              // текущая строка
   reg[2:0] fontcol;          // столбец шрифта
   reg[4:0] fontrow;          // строка шрифта
   reg[12:0] char_adr;       // адрес текущего знакоместа в видеопамяти
   reg[12:0] row_start_adr;   // адрес начала текущей строки в виедопамяти
   reg[3:0] cursor_match;         // флаг наличия курсора в текущей позиции
   reg[7:0] char_evn;             // четный символ
   reg[7:0] char_odd;             // нечетный символ
   reg[14:0] font_adr;            // адрес в шрифтовой памяти
   wire pixel;                    // выход данных шрифтовой памяти
   reg vram_a0_selector;  // признак четного-нечетного знакоместа
	reg vga_out;           // регистр видеосигнала -состояние теущего пикселя (0 - откл, 1 - вкл)
	wire cursor_pixel;     // признак вывода курсорных пикселей
	wire cursor_pixel_d;   // тот же сигнал с задержкой в 1 пиксель
   wire cursor_field;     // признак вывода строк, на которых разрешено отображение курсора
   reg [1:0] flashflag;   // признак вывода данного символа мерцающим	
	
	// ограничитель счетчика строк для одного знакоместа в зависимости от числа отображаемых строк
	wire[5:0] fontrowlimit;        
	assign fontrowlimit = (lmode == 0)? 5'd17:5'd11;
	
	// Селектор цветов выводимого видеосигнала
   assign vgab = ((char_adr < 13'd159) && (char_adr> 13'd70))  ? vga_out:1'b0;  // синий - часы и разделительная черта
   assign vgar = ((row_start_adr == 13'b0) || cursor_pixel_d)? vga_out:1'b0;      // красный - служебная строка и курсор 
	assign vgag = (row_start_adr > 13'd159)? vga_out:1'b0;                         // зеленый - все строки начиная с 2
   // признак наличия курсора в данном пикселе  
	assign cursor_field = (fontrow[3:1] == 3'b101) | cursor_type; // для строк 10-11 или все знакоместо
	assign cursor_pixel= cursor_match[2] && cursor_field;
	assign cursor_pixel_d= cursor_match[3] && cursor_field;
	
   //************************************
   //* ROM знакогенератора с шрифтами 
   //************************************
   fontrom fontrom0 (
      .address(font_adr), 
      .clock(vgaclk), 
      .q(pixel)
   ); 

   //**********************************************
	// Генератор основной пиксельной частоты 25 Мгц
   //**********************************************	
   always @(posedge clk50mhz) begin
      if (wb_rst_i == 1'b1) vgaclk <= 1'b0 ;   // после сброса начинаем с 0
      else  vgaclk <= ~vgaclk ;   // инвертируем сигнал каждый перепад 50 Мгц
   end 

	//**********************************************
	//* Связь с шиной
	//**********************************************
	wire bus_strobe = wb_cyc_i & wb_stb_i;         // строб цикла шины
	wire bus_read_req = bus_strobe & ~wb_we_i;     // запрос чтения
	wire bus_write_req = bus_strobe & wb_we_i;     // запрос записи

   // формирователь ответа на цикл шины	
	wire reply=wb_cyc_i & wb_stb_i & ~wb_ack_o;
	
	// Сигнал ответа 
	always @(posedge wb_clk_i or posedge wb_rst_i)
     if (wb_rst_i == 1) wb_ack_o <= 0;
	  else wb_ack_o <= reply;

	// обработка шинных транзакций  
   always @(posedge wb_clk_i)  begin
	   
	   // Чтение данных из видеопамяти
      if (bus_read_req == 1'b1) begin
        wb_dat_o[7:0] <= vram_even[wb_adr_i[12:1]] ; 
        wb_dat_o[15:8] <= vram_odd[wb_adr_i[12:1]] ;
	   end
      // запись данных в видеопамять	
      if (bus_write_req == 1'b1)  begin
		   // запись четных байтов 
         if (wb_sel_i[0] == 1'b1) vram_even[wb_adr_i[12:1]] <= wb_dat_i[7:0] ; 
		   // запись нечетных байтов
         if (wb_sel_i[1] == 1'b1) vram_odd[wb_adr_i[12:1]] <= wb_dat_i[15:8] ; 
      end  
   end 

	//********************************************
	//* Формирователь видеосигнала  640*480
	//********************************************
   always @(posedge vgaclk)  begin
	   // Сброс видеоформирователя
      if (wb_rst_i == 1'b1)  begin
         col <= 0 ; 
         row <= 0 ; 
         row_start_adr <= 13'b0000000000000 ; 
         fontrow <= 5'b00000 ; 
         vga_hsync <= 1'b1 ; 
         vga_vsync <= 1'b1 ; 
         vga_out <= 1'b0 ; 
			flashflag <= 2'b11;
      end
		
		//**************************************
		// попиксельная обработка
		//**************************************
      else  begin
		   // Счетчик колонок - строчная развертка, 800 точек в строке (640  видимых и 160 служебных)
			//----------------------------------------------------------------------------------------------
         if (col < 11'd799) col <= col + 1'b1 ; // переход на следующий пиксель

         //**************************************
			// переход на новую строку
         //**************************************
         else begin
            col <= 0 ; // колонка 0
				// счетчик колонок знакоместа - 8 точек шрифта, остальное - межстрочный интервал
            if (fontrow < fontrowlimit) fontrow <= fontrow + 1'b1 ; 
            else begin
				   // переход на новое знакоместо
               fontrow <= 5'b00000 ; 
               row_start_adr <= row_start_adr + 7'd80 ; // адрес в видеобуфере+80 - следующая строка (строки по 80 байт)
            end 
				
				// Счетчик строк - кадровая развертка, 524 строки (480 видимых и 44 служебных)
				//--------------------------------------------------------------------------------
            if (row < 10'd523) begin
				   // вывод строк видимой части кадра
               row <= row + 1'b1 ; // следующая строка
               if (row >= 10'd479) begin
					   // конец видимой части кадра
                  row_start_adr <= 13'b0000000000000 ; 
                  fontrow <= 5'b00000 ; 
               end 
            end
				
    		   // Переход на новый кадр	
            else  begin
               row <= 10'd0 ; // строка 0
               row_start_adr <= 13'b0000000000000 ; // начало строки в видеобуфере
               fontrow <= 5'b00000 ;            // первая точка шрифта строки
            end 
         end

			//********************************************
		   // Строчная синхронизация, начало строки
			//********************************************
			// столбцы 00-95
         vga_out <= 1'b0 ;   // отключаем видеосигнал
         if (col < 11'd96) vga_hsync <= 1'b0 ; // первые 95 столбцов - строчный синхроимпульс

			//*************************************************
		   // Гашение сигнала после строчного синхроимпульса
			//*************************************************
         // столбцы 96-140			
         else if (col < 11'd141)  begin
            vga_hsync <= 1'b1 ; // снимаем строчный синхроимпульс
            fontcol <= 3'b000 ;      // подготавливаем счетчик колонок шрифта 
            char_adr <= row_start_adr ; // адрес текущего символа равен адресу начала строки
         end
			
			//********************************************
		   // Формирователь видимой части строки
			//********************************************
			// столбцы 141-783
         else if (col < 11'd784)  begin
			   // строка текущего символа отрисована - переход к следующему символу
            if (fontcol == 3'b110)  char_adr <= char_adr + 1'b1 ; 
				
				// последовательный перебор всех точек шрифта текущего символа - от 0 до 7
            fontcol <= fontcol + 1'b1 ; 
				
				// 144 колонка - гашение видеосигнала по обратному ходу
            if (col < 11'd144)    vga_out <= 1'b0 ;  

			   // запись регистра видеовыхода
            else 	if (fontrow < 4'd12) begin
				  // пиксели,занимаемые курсором, имеют инверсию видеосигнала
              if (cursor_pixel) vga_out <= ~pixel; 
				  // формирование обычных пикселей с учетом флага мерцания
  				  else   vga_out <= pixel & (flash | flashflag[1]) ; 
				end  
				// межстрочные промежутки
				else vga_out <= 1'b0;  
         end

			//********************************
			// обработка курсора
			//********************************
         if ((char_adr == cursor) & cursor_on)  cursor_match <= {cursor_match[2:0], 1'b1} ; // вводим признак курсора в сдвиговый регистр
         else                                   cursor_match <= {cursor_match[2:0], 1'b0} ; // курсора нет - начинаем заполнять регистр нулями
       
			//***************************************************
		   // формирователь адреса пикселя в массиве шрифтов	
			//***************************************************
         // определение четных-нечетных байтов			
         if ((char_adr[0]) == 1'b0)   vram_a0_selector <= 1'b0 ; // четные знакосимволы
         else                         vram_a0_selector <= 1'b1 ; // нечетные
         // выборка четного и нечетного байта из видеопамяти
         char_evn <= vram_even[char_adr[12:1]] ; // четный теущий символ
         char_odd <= vram_odd[char_adr[12:1]] ; // нечетный текущий символ
         // формирование адреса текущей точки в массиве шрифтов
         if (vram_a0_selector == 1'b0)  font_adr <= ({fontrow[3:0], 11'b00000000000}) | ({fontcol, 8'b00000000}) | char_evn ; // четные символы
         else                           font_adr <= ({fontrow[3:0], 11'b00000000000}) | ({fontcol, 8'b00000000}) | char_odd ; // нечетные символы

			//********************************************
         //*  Формирователь флага мерцания символов
			//********************************************
	      // Флаг формируется для символов с кодами 00-1F		
         if ((vram_a0_selector == 1'b0) && (char_evn[7:5] == 3'b000) ||  // для четных символов
			    (vram_a0_selector == 1'b1) && (char_odd[7:5] == 3'b000))    // для нечетных символов
				   flashflag[0] <= 1'b0;  // флаг поднят (0)
         else  flashflag[0] <= 1'b1;  // для остальных флаг опущен (1)
			flashflag[1] <= flashflag[0]; // задержка флага на 1 пиксель
			
			//***************************************************************
         //*  Кадровая синхронизация
			//***************************************************************
         if (row > 10'd479)  vga_out <= 1'b0 ;  // на строках выше 479 видеосигнала нет 
			// строки 480-489 - гашение перед синхроимпульсом (front porch)
			// строка 490 - кадровый синхроимпульс
   		if (row == 10'd490) vga_vsync <= 1'b0 ;  
         else                vga_vsync <= 1'b1 ; 
         // оставшиеся 34 строки - гашение после синхроимпульса (back porch)  - обратный ход кадровой развертки
			
			
      end  
   end 
endmodule
